module add(input [15:0] a,b, output reg [15:0] result);

	always@(*)

	beging 
		result = a + b; 
	end 

endmodule