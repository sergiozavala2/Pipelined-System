`include "alu.v"

module alu_tb;


alu utt(a, b, function, out, r15);

initial 
begin 

$monitor()

end 

initial
begin

//signed addition 
#10 

//signed subtraction 

//signed multiplication 

//signed division 
